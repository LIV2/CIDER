localparam  Z2_IDLE  = 2'd0,
            Z2_START = 2'd1,
            Z2_DATA  = 2'd2,
            Z2_END   = 2'd3;